`define FNADD  0
`define FNSL	1
`define FNLR	2
`define FNSEQ	2
`define FNSC   3
`define FNSNE	3
`define FNXOR	4
`define FNSR	5
`define FNOR	6
`define FNAND	7
`define FNSUB	10
`define FNSRA	11
`define FNSLT	12
`define FNSGE	13
`define FNSLTU	14
`define FNSGEU	15

`define FNSWAP 1 
`define FMINU	10
`define FMIN	11
`define FMAXU  12
`define FMAX	13

`define FNRAND	8
